module testactor

pub fn (mut actor Testactor) transform_base_object(base_object BaseObject) ! {
	// some custom function on base object
}
