module testactor

pub struct AnotherObject {
	text   string
	number int @[index]
}
