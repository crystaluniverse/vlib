module main

import os
import time

pub struct App {
pub:
	secret_key string = '1234'
}

pub fn main() {
	// mut app := App{
	// }
	println('Hello V')
	time.sleep(1 * time.hour)
	println('Goodbye V')
}
