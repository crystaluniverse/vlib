module openrouter

// https://openrouter.ai/docs/models
// todo: see also /root/code/github/freeflowuniverse/crystallib/crystallib/clients/openai/models.v
