module canva

// cmd:='curl -X GET "https://api.canva.com/v1/designs/DESIGN_ID/download" -H "Authorization: Bearer YOUR_ACCESS_TOKEN" -H "Content-Type: application/json"''
